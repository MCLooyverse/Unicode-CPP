Lu|kLetterUppercase
Ll|kLetterLowercase
Lt|kLetterTitlecase
Lm|kLetterModifier
Lo|kLetterOther
Mn|kMarkNonspacing
Mc|kMarkSpacingCombining
Me|kMarkEnclosing
Nd|kNumberDecimalDigit
Nl|kNumberLetter
No|kNumberOther
Pc|kPunctuationConnector
Pd|kPunctuationDash
Ps|kPunctuationOpen
Pe|kPunctuationClose
Pi|kPunctuationInitialQuote
Pf|kPunctuationFinalQuote
Po|kPunctuationOther
Sm|kSymbolMath
Sc|kSymbolCurrency
Sk|kSymbolModifier
So|kSymbolOther
Zs|kSeparatorSpace
Zl|kSeparatorLine
Zp|kSeparatorParagraph
Cc|kOtherControl
Cf|kOtherFormat
Cs|kOtherSurrogate
Co|kOtherPrivateUse
Cn|kOtherNotAssigned
